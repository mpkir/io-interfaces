

module a_black_box (
	input [ 1:0]  ctrl,
	inout [23:0]  iopad_a,
	inout [23:0]  iopad_b
);

// logic internal to black box not shown

endmodule

